//Debouncer

module debounce(input logic clk, signal_in output logic signal_out);


endmodule